`include "float_adder.v"

module test_float_adder;
    reg clk = 1;
    always #5 clk = ~clk;
    reg [31:0] a, b;
    wire [31:0] c;
    wire [2:0] state;
    reg rst;
    reg [31:0] a_array [0:99];
    reg [31:0] b_array [0:99];
    reg [31:0] c_array [0:99];
    FAdd float_adder(
        .clk(clk),
        .rst(rst),
        .a(a),
        .b(b),
        .c(c),
        .state(state)
    );
    integer i;
    integer j;
    initial begin
    a_array[0] = 32'b10111111010101110001011010001011;
    b_array[0] = 32'b00111111010010000111100100110001;
    c_array[0] = 32'b10111101011010011101010110100000;
    a_array[1] = 32'b00111111011010010110000110111001;
    b_array[1] = 32'b10111110101010111010001001010001;
    c_array[1] = 32'b00111111000100111001000010010000;
    a_array[2] = 32'b00111110100011100011100001111101;
    b_array[2] = 32'b00111110111101000110110101100011;
    c_array[2] = 32'b00111111010000010101001011110000;
    a_array[3] = 32'b00111110101110101100010100001000;
    b_array[3] = 32'b10111111011100111100010101010100;
    c_array[3] = 32'b10111111000101100110001011010000;
    a_array[4] = 32'b10111111001000101011111000000001;
    b_array[4] = 32'b10111110000100010000000001000011;
    c_array[4] = 32'b10111111010001101111111000010010;
    a_array[5] = 32'b10111100100001011000100011000111;
    b_array[5] = 32'b00111110000011001000011001101111;
    c_array[5] = 32'b00111101111101111010101010101100;
    a_array[6] = 32'b10111110001000000111000001111100;
    b_array[6] = 32'b00111110000001001110011111001001;
    c_array[6] = 32'b10111100110111000100010110011000;
    a_array[7] = 32'b00111111011111111011100110000100;
    b_array[7] = 32'b10111111000000110100111110001010;
    c_array[7] = 32'b00111110111110001101001111110100;
    a_array[8] = 32'b10111111000111001101010111110111;
    b_array[8] = 32'b00111111001000110011011010100000;
    c_array[8] = 32'b00111100110011000001010100100000;
    a_array[9] = 32'b10111110111111001011011011101001;
    b_array[9] = 32'b10111110100101011100010011000011;
    c_array[9] = 32'b10111111010010010011110111010110;
    a_array[10] = 32'b00111111000001101101100011000010;
    b_array[10] = 32'b00111110110011001110101011000100;
    c_array[10] = 32'b00111111011011010100111000100100;
    a_array[11] = 32'b00111110100100010000111010100001;
    b_array[11] = 32'b10111111010011101100011100001001;
    c_array[11] = 32'b10111111000001100011111110111000;
    a_array[12] = 32'b10111101100011101101101111011011;
    b_array[12] = 32'b10111111000001101010011110100010;
    c_array[12] = 32'b10111111000110001000001100011101;
    a_array[13] = 32'b10111110010001001101001110110101;
    b_array[13] = 32'b00111111011000111110011001001001;
    c_array[13] = 32'b00111111001100101011000101011100;
    a_array[14] = 32'b10111101100000110110110001000001;
    b_array[14] = 32'b00111110111010100101011111100010;
    c_array[14] = 32'b00111110110010010111110011010010;
    a_array[15] = 32'b00111110011100111111111110101001;
    b_array[15] = 32'b00111111011001101111011100011100;
    c_array[15] = 32'b00111111100100011111101110000011;
    a_array[16] = 32'b00111110100010001000100001101010;
    b_array[16] = 32'b00111110110000000001101100100001;
    c_array[16] = 32'b00111111001001000101000111000110;
    a_array[17] = 32'b00111111000000110011010110000101;
    b_array[17] = 32'b00111111000010000001011101011100;
    c_array[17] = 32'b00111111100001011010011001110000;
    a_array[18] = 32'b00111110111000000001001000001001;
    b_array[18] = 32'b00111111011011100100100110001101;
    c_array[18] = 32'b00111111101011110010100101001001;
    a_array[19] = 32'b10111110100100011000111011101000;
    b_array[19] = 32'b10111111001000111101010110100111;
    c_array[19] = 32'b10111111011011001001110100011011;
    a_array[20] = 32'b10111111001100000001011110101111;
    b_array[20] = 32'b10111110111000010101010101100001;
    c_array[20] = 32'b10111111100100000110000100110000;
    a_array[21] = 32'b10111111010101000100011010000110;
    b_array[21] = 32'b00111110011010100111011010100010;
    c_array[21] = 32'b10111111000110011010100011011110;
    a_array[22] = 32'b00111110101100110110001001101001;
    b_array[22] = 32'b10111111011101001101101100011010;
    c_array[22] = 32'b10111111000110110010100111100110;
    a_array[23] = 32'b10111111001010000100010100010100;
    b_array[23] = 32'b10111110111000010000110111111111;
    c_array[23] = 32'b10111111100011000110011000001010;
    a_array[24] = 32'b10111110110010111111111111100100;
    b_array[24] = 32'b00111111001011110010100011110010;
    c_array[24] = 32'b00111110100100100101001000000000;
    a_array[25] = 32'b10111110111101110000100100000100;
    b_array[25] = 32'b10111111011100110100001110111101;
    c_array[25] = 32'b10111111101101110110010000100000;
    a_array[26] = 32'b00111110000101110011010000110000;
    b_array[26] = 32'b10111111001001000001110111011100;
    c_array[26] = 32'b10111110111111001010000110100000;
    a_array[27] = 32'b10111111000111101001110111100000;
    b_array[27] = 32'b10111111010010010011011101101111;
    c_array[27] = 32'b10111111101100111110101010101000;
    a_array[28] = 32'b10111110111001001110000110010110;
    b_array[28] = 32'b00111110010000000000100010101110;
    c_array[28] = 32'b10111110100001001101110100111111;
    a_array[29] = 32'b00111111000011100111001100011001;
    b_array[29] = 32'b00111110001011011010110101111011;
    c_array[29] = 32'b00111111001110011101111001111000;
    a_array[30] = 32'b00111101110100110100101101101010;
    b_array[30] = 32'b00111110111111011010101011011000;
    c_array[30] = 32'b00111111000110010011111011011001;
    a_array[31] = 32'b00111111011111000001100010101111;
    b_array[31] = 32'b00111111001011110011011111001010;
    c_array[31] = 32'b00111111110101011010100000111100;
    a_array[32] = 32'b00111111001111111111000011111100;
    b_array[32] = 32'b10111110100101101001110000110000;
    c_array[32] = 32'b00111110111010010100010111001000;
    a_array[33] = 32'b00111111000101011010000100001010;
    b_array[33] = 32'b00111110000111000000110000010010;
    c_array[33] = 32'b00111111001111001010010000001110;
    a_array[34] = 32'b00111110000000000111110001111110;
    b_array[34] = 32'b10111110001010000000101001010110;
    c_array[34] = 32'b10111101000111100011011101100000;
    a_array[35] = 32'b00111101100110001010001100010100;
    b_array[35] = 32'b00111101010101110010100011101100;
    c_array[35] = 32'b00111110000000100001101111000101;
    a_array[36] = 32'b00111110001101000111000010010001;
    b_array[36] = 32'b10111111010011000011110001111110;
    c_array[36] = 32'b10111111000111110010000001011010;
    a_array[37] = 32'b00111111001010000001010010001110;
    b_array[37] = 32'b00111111001000111011001110001011;
    c_array[37] = 32'b00111111101001011110010000001100;
    a_array[38] = 32'b00111101101111110111001010110001;
    b_array[38] = 32'b00111111000001010010110001111101;
    c_array[38] = 32'b00111111000111010001101011010011;
    a_array[39] = 32'b00111101100011110010101100010110;
    b_array[39] = 32'b00111110111011000011111101001110;
    c_array[39] = 32'b00111111000010000000010100001010;
    a_array[40] = 32'b10111111000100101100010100000010;
    b_array[40] = 32'b10111101010101001011110111001100;
    c_array[40] = 32'b10111111001000000001000011011111;
    a_array[41] = 32'b10111111011111111111111110010100;
    b_array[41] = 32'b10111111011000111101010000100010;
    c_array[41] = 32'b10111111111100011110100111011011;
    a_array[42] = 32'b10111111011111110110111111000001;
    b_array[42] = 32'b10111111010111101101101110110011;
    c_array[42] = 32'b10111111111011110010010110111010;
    a_array[43] = 32'b10111011100010000101111000011011;
    b_array[43] = 32'b00111111000110000000100101010001;
    c_array[43] = 32'b00111111000101101111100010010101;
    a_array[44] = 32'b00111110001001110000101111110010;
    b_array[44] = 32'b10111111011010011011110000011110;
    c_array[44] = 32'b10111111001111111111100100100010;
    a_array[45] = 32'b00111110101101111101101101011001;
    b_array[45] = 32'b10111111000101000101010110000110;
    c_array[45] = 32'b10111110011000011001111101100110;
    a_array[46] = 32'b00111111001011111111100010011111;
    b_array[46] = 32'b00111111000001111110001100001000;
    c_array[46] = 32'b00111111100110111110110111010100;
    a_array[47] = 32'b00111110100110111100110010010011;
    b_array[47] = 32'b00111111000100111011010001100001;
    c_array[47] = 32'b00111111011000011001101010101010;
    a_array[48] = 32'b00111111001111110111000001101110;
    b_array[48] = 32'b10111101000100010001010110000011;
    c_array[48] = 32'b00111111001101100101111100010110;
    a_array[49] = 32'b00111111010101010100111100011111;
    b_array[49] = 32'b00111111010111111000111010110110;
    c_array[49] = 32'b00111111110110100110111011101010;
    a_array[50] = 32'b01111101010111100001100011111000;
    b_array[50] = 32'b11110011101000011000001000011011;
    c_array[50] = 32'b01111101010111100001100011100100;
    a_array[51] = 32'b01010101010111000101010110110101;
    b_array[51] = 32'b00010100111111001110011101001110;
    c_array[51] = 32'b01010101010111000101010110110101;
    a_array[52] = 32'b01110001110010010001001010011000;
    b_array[52] = 32'b01010011001010011001100100111000;
    c_array[52] = 32'b01110001110010010001001010011000;
    a_array[53] = 32'b11010000100100101100101001111001;
    b_array[53] = 32'b01011001101011011110101000111101;
    c_array[53] = 32'b01011001101011011110101000011000;
    a_array[54] = 32'b10101010000101010101110110111100;
    b_array[54] = 32'b10001001011111100001101101001110;
    c_array[54] = 32'b10101010000101010101110110111100;
    a_array[55] = 32'b10011100101000001100010111111010;
    b_array[55] = 32'b11000001010111100010100001101100;
    c_array[55] = 32'b11000001010111100010100001101100;
    a_array[56] = 32'b00100011110110000110101010101100;
    b_array[56] = 32'b11011100000100001111111000100001;
    c_array[56] = 32'b11011100000100001111111000100001;
    a_array[57] = 32'b00111100010110011001000110101010;
    b_array[57] = 32'b01111000110111110110101001010101;
    c_array[57] = 32'b01111000110111110110101001010101;
    a_array[58] = 32'b00101011000011011000110110111110;
    b_array[58] = 32'b10110111100111100010000110110101;
    c_array[58] = 32'b10110111100111100010000110110101;
    a_array[59] = 32'b00101100001001110001011100111011;
    b_array[59] = 32'b11101010101001111011011101011100;
    c_array[59] = 32'b11101010101001111011011101011100;
    a_array[60] = 32'b01010110011101011111111100110110;
    b_array[60] = 32'b10111101101100000001001010110011;
    c_array[60] = 32'b01010110011101011111111100110110;
    a_array[61] = 32'b01011011001001011010110011100010;
    b_array[61] = 32'b01001111100101111110001111100100;
    c_array[61] = 32'b01011011001001011010110011100011;
    a_array[62] = 32'b00110100111111010110101101001111;
    b_array[62] = 32'b11010110010000111000110100010101;
    c_array[62] = 32'b11010110010000111000110100010101;
    a_array[63] = 32'b00101100011011100100101011111101;
    b_array[63] = 32'b11001101111101110010111001001110;
    c_array[63] = 32'b11001101111101110010111001001110;
    a_array[64] = 32'b01011101100010001000101000001000;
    b_array[64] = 32'b01011110110001101010111111010100;
    c_array[64] = 32'b01011110111010001101001001010110;
    a_array[65] = 32'b11110101111000001000010110001010;
    b_array[65] = 32'b01010011100110011100011001010100;
    c_array[65] = 32'b11110101111000001000010110001010;
    a_array[66] = 32'b01000100001001110000011010011010;
    b_array[66] = 32'b10100001010101111111011010111100;
    c_array[66] = 32'b01000100001001110000011010011010;
    a_array[67] = 32'b01010111110100101111000100001110;
    b_array[67] = 32'b00001110001111100100011110101000;
    c_array[67] = 32'b01010111110100101111000100001110;
    a_array[68] = 32'b11001001110100001111111010101100;
    b_array[68] = 32'b01010101010100011011100111110011;
    c_array[68] = 32'b01010101010100011011100111110001;
    a_array[69] = 32'b11100011010011000101011101001100;
    b_array[69] = 32'b10101010001100011011011000101101;
    c_array[69] = 32'b11100011010011000101011101001100;
    a_array[70] = 32'b01111101111111111001110100001001;
    b_array[70] = 32'b01101001111001111111001111100101;
    c_array[70] = 32'b01111101111111111001110100001001;
    a_array[71] = 32'b10011000000101101111100011000100;
    b_array[71] = 32'b11111010101101001001110110101111;
    c_array[71] = 32'b11111010101101001001110110101111;
    a_array[72] = 32'b01100001111001110100111010100011;
    b_array[72] = 32'b10001111100000011001111001111111;
    c_array[72] = 32'b01100001111001110100111010100011;
    a_array[73] = 32'b00110001001000010110011110101101;
    b_array[73] = 32'b11111000101101011110011101110110;
    c_array[73] = 32'b11111000101101011110011101110110;
    a_array[74] = 32'b01101110010100110100110011011110;
    b_array[74] = 32'b01100101100101101000110000011100;
    c_array[74] = 32'b01101110010100110100110100101001;
    a_array[75] = 32'b00100110000011011000110001001010;
    b_array[75] = 32'b01110100011011110010111000110000;
    c_array[75] = 32'b01110100011011110010111000110000;
    a_array[76] = 32'b10111111110000110010111000100000;
    b_array[76] = 32'b00010100110101010011011010000101;
    c_array[76] = 32'b10111111110000110010111000100000;
    a_array[77] = 32'b01101110101010101000010111111011;
    b_array[77] = 32'b00111011010110010100100000000111;
    c_array[77] = 32'b01101110101010101000010111111011;
    a_array[78] = 32'b00111111011111000010111111110100;
    b_array[78] = 32'b10010111000110000000101100001011;
    c_array[78] = 32'b00111111011111000010111111110100;
    a_array[79] = 32'b01011101001000000101111000100000;
    b_array[79] = 32'b11001101001100101010101110000110;
    c_array[79] = 32'b01011101001000000101111000100000;
    a_array[80] = 32'b11101011010001111111011000111110;
    b_array[80] = 32'b00010110110011111000000011110001;
    c_array[80] = 32'b11101011010001111111011000111110;
    a_array[81] = 32'b10111111110011111010111011011001;
    b_array[81] = 32'b10010001101100011100110000110011;
    c_array[81] = 32'b10111111110011111010111011011001;
    a_array[82] = 32'b00101001100100110100011010011001;
    b_array[82] = 32'b11110100010010010011100110100011;
    c_array[82] = 32'b11110100010010010011100110100011;
    a_array[83] = 32'b11101011000111010010110000010100;
    b_array[83] = 32'b00111111011111110101110111011001;
    c_array[83] = 32'b11101011000111010010110000010100;
    a_array[84] = 32'b00110010011110010100111111110111;
    b_array[84] = 32'b01001101111011111101111110100000;
    c_array[84] = 32'b01001101111011111101111110100000;
    a_array[85] = 32'b00010011010110111000000100010000;
    b_array[85] = 32'b10001101110011011111100011110110;
    c_array[85] = 32'b00010011010110110110011101010001;
    a_array[86] = 32'b10101110100010100110001110010100;
    b_array[86] = 32'b00101010011010101101100110111110;
    c_array[86] = 32'b10101110100010011110111000100111;
    a_array[87] = 32'b00110110101100101010110010111100;
    b_array[87] = 32'b01001010101100100110111001111000;
    c_array[87] = 32'b01001010101100100110111001111000;
    a_array[88] = 32'b11010100010100011100111101001001;
    b_array[88] = 32'b10111110011001000000000011100110;
    c_array[88] = 32'b11010100010100011100111101001001;
    a_array[89] = 32'b01110001000001110101011111010000;
    b_array[89] = 32'b11000010010001000111100111011010;
    c_array[89] = 32'b01110001000001110101011111010000;
    a_array[90] = 32'b01000111010111100010010101101010;
    b_array[90] = 32'b01101010001110110111000101001100;
    c_array[90] = 32'b01101010001110110111000101001100;
    a_array[91] = 32'b10011111010001100001101101010001;
    b_array[91] = 32'b01011101010110111010101110110011;
    c_array[91] = 32'b01011101010110111010101110110011;
    a_array[92] = 32'b11111110000011110110001110000100;
    b_array[92] = 32'b01110010111000110100000100111010;
    c_array[92] = 32'b11111110000011110110001110000010;
    a_array[93] = 32'b10110100100101001011001011111011;
    b_array[93] = 32'b01100100010000101001010110011001;
    c_array[93] = 32'b01100100010000101001010110011001;
    a_array[94] = 32'b10100101100101110011111000110010;
    b_array[94] = 32'b01101110110010011101100001000100;
    c_array[94] = 32'b01101110110010011101100001000100;
    a_array[95] = 32'b00000110010010101111010010011011;
    b_array[95] = 32'b11111110010001001000110111101001;
    c_array[95] = 32'b11111110010001001000110111101001;
    a_array[96] = 32'b10011010111111100011011000100101;
    b_array[96] = 32'b11101110101111100100001000001000;
    c_array[96] = 32'b11101110101111100100001000001000;
    a_array[97] = 32'b00001100101111100101101111101001;
    b_array[97] = 32'b10001100101111100101101111101001;
    c_array[97] = 32'b00000000000000000000000000000000;
    a_array[98] = 32'b00000000000000000000000000000000;
    b_array[98] = 32'b10000000000000000000000000000000;
    c_array[98] = 32'b00000000000000000000000000000000;
    a_array[99] = 32'b11111111100000000000000000000000;
    b_array[99] = 32'b01111111100000000000000000000000;
    c_array[99] = 32'b01111111100000000000000000000001;
        #5;
        for (i = 0; i < 100; i = i + 1) begin
            rst = 0;
            #10;
            rst = 1;
            a = a_array[i];
            b = b_array[i];
            for (j = 0; j < 300; j = j + 1) begin // it takes at most about 255 + 32 cycles to finish the calculation
//                $display("state: %d, c: %b", state, c);
                #10;
            end
            if (c !== c_array[i] && !(c === 32'b01111111100000000000000000000001 && c_array[i][30:23] === 8'b11111111 && c_array[i][22:0] !== 23'b0)) begin
                 $display("Wrong Answer! i: %d, a: %b, b: %b, output: %b, expected: %b", i, a, b, c, c_array[i]);
                 $fatal;
            end
        end
		$display("Congratulations! You have passed all of the tests.");
		$finish;
    end
endmodule