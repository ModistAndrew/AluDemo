`include "float_adder.v"

module test_float_adder;
    reg clk = 1;
    always #5 clk = ~clk;
    reg [31:0] a, b;
    wire [31:0] c;
    wire [2:0] state;
    reg rst;
    reg [31:0] a_array [0:99];
    reg [31:0] b_array [0:99];
    reg [31:0] c_array [0:99];
    FAdd float_adder(
        .clk(clk),
        .rst(rst),
        .a(a),
        .b(b),
        .c(c),
        .state(state)
    );
    integer i;
    integer j;
    initial begin
        #5;
        a_array[0] = 32'b0;
        b_array[0] = 32'b0;
        c_array[0] = 32'b0;
        a_array[1] = 32'b00111111010010000111100100110001;
        b_array[1] = 32'b00111111010011000110011010010001;
        c_array[1] = 32'b00111111110010100110111111100001;
        a_array[2] = 32'b00111111011010010110000110111001;
        b_array[2] = 32'b00111110010010100100101011101000;
        c_array[2] = 32'b00111111100011011111101000111010;
        a_array[3] = 32'b00111110101010111010001001010001;
        b_array[3] = 32'b00111111010001001010101010110010;
        c_array[3] = 32'b00111111100011010011110111101101;
        a_array[4] = 32'b00111110100011100011100001111101;
        b_array[4] = 32'b00111111000011011101000011111010;
        c_array[4] = 32'b00111111010101001110110100111000;
        a_array[5] = 32'b00111110111101000110110101100011;
        b_array[5] = 32'b00111111001000001111110110101111;
        c_array[5] = 32'b00111111100011011001101000110000;
        a_array[6] = 32'b00111110101110101100010100001000;
        b_array[6] = 32'b00111111000000110110111000111110;
        c_array[6] = 32'b00111111011000001101000011000010;
        a_array[7] = 32'b00111111011100111100010101010100;
        b_array[7] = 32'b00111111011010101000101111000011;
        c_array[7] = 32'b00111111111011110010100010001100;
        a_array[8] = 32'b00111111001000101011111000000001;
        b_array[8] = 32'b00111111001101111010000011000110;
        c_array[8] = 32'b00111111101011010010111101100100;
        a_array[9] = 32'b00111110000100010000000001000011;
        b_array[9] = 32'b00111111000110110110001001010000;
        c_array[9] = 32'b00111111001111111010001001100001;
        a_array[10] = 32'b00111100100001011000100011000111;
        b_array[10] = 32'b00111110011110001011011101001111;
        c_array[10] = 32'b00111110100001001011010000110100;
        a_array[11] = 32'b00111110000011001000011001101111;
        b_array[11] = 32'b00111111010011011101111010000111;
        c_array[11] = 32'b00111111011100010000000000100011;
        a_array[12] = 32'b00111110001000000111000001111100;
        b_array[12] = 32'b00111110110011010100100010010101;
        c_array[12] = 32'b00111111000011101100000001101010;
        a_array[13] = 32'b00111110000001001110011111001001;
        b_array[13] = 32'b00111101110111101101011100100110;
        c_array[13] = 32'b00111110011101000101001101011100;
        a_array[14] = 32'b00111111011111111011100110000100;
        b_array[14] = 32'b00111110010111110111111010111101;
        c_array[14] = 32'b00111111100110111100110010011010;
        a_array[15] = 32'b00111111000000110100111110001010;
        b_array[15] = 32'b00111111010101101101000000001111;
        c_array[15] = 32'b00111111101011010000111111001100;
        a_array[16] = 32'b00111111000111001101010111110111;
        b_array[16] = 32'b00111110100101111001000101110101;
        c_array[16] = 32'b00111111011010001001111010110010;
        a_array[17] = 32'b00111111001000110011011010100000;
        b_array[17] = 32'b00111111000001100011011110101111;
        c_array[17] = 32'b00111111100101001011011100101000;
        a_array[18] = 32'b00111110111111001011011011101001;
        b_array[18] = 32'b00111111011110010000011111001001;
        c_array[18] = 32'b00111111101110111011000110011111;
        a_array[19] = 32'b00111110100101011100010011000011;
        b_array[19] = 32'b00111111010001010111011110110011;
        c_array[19] = 32'b00111111100010000010110100001010;
        a_array[20] = 32'b00111111000001101101100011000010;
        b_array[20] = 32'b00111111010001010001100100010011;
        c_array[20] = 32'b00111111101001011111100011101010;
        a_array[21] = 32'b00111110110011001110101011000100;
        b_array[21] = 32'b00111111011001000011101101000110;
        c_array[21] = 32'b00111111101001010101100001010100;
        a_array[22] = 32'b00111110100100010000111010100001;
        b_array[22] = 32'b00111110101101000111010101101100;
        c_array[22] = 32'b00111111001000101100001000000110;
        a_array[23] = 32'b00111111010011101100011100001001;
        b_array[23] = 32'b00111111011010110100010101010010;
        c_array[23] = 32'b00111111110111010000011000101110;
        a_array[24] = 32'b00111101100011101101101111011011;
        b_array[24] = 32'b00111111011100110000011100011001;
        c_array[24] = 32'b00111111100000100111000101001010;
        a_array[25] = 32'b00111111000001101010011110100010;
        b_array[25] = 32'b00111101101100000011111000001100;
        c_array[25] = 32'b00111111000111001010111101100100;
        a_array[26] = 32'b00111110010001001101001110110101;
        b_array[26] = 32'b00111111001010011100100100111101;
        c_array[26] = 32'b00111111010110101111111000101010;
        a_array[27] = 32'b00111111011000111110011001001001;
        b_array[27] = 32'b00111110101100101010001000011000;
        c_array[27] = 32'b00111111100111101001101110101010;
        a_array[28] = 32'b00111101100000110110110001000001;
        b_array[28] = 32'b00111100101001000000011101100000;
        c_array[28] = 32'b00111101101011000110111000011001;
        a_array[29] = 32'b00111110111010100101011111100010;
        b_array[29] = 32'b00111101100000010011100001100100;
        c_array[29] = 32'b00111111000001010101001011111110;
        a_array[30] = 32'b00111110011100111111111110101001;
        b_array[30] = 32'b00111111011110000111101101111010;
        c_array[30] = 32'b00111111100110101011110110110010;
        a_array[31] = 32'b00111111011001101111011100011100;
        b_array[31] = 32'b00111111010110011101010111100001;
        c_array[31] = 32'b00111111111000000110011001111110;
        a_array[32] = 32'b00111110100010001000100001101010;
        b_array[32] = 32'b00111111000010100010110110111100;
        c_array[32] = 32'b00111111010011100111000111110001;
        a_array[33] = 32'b00111110110000000001101100100001;
        b_array[33] = 32'b00111111010000101001111110101001;
        c_array[33] = 32'b00111111100100010101011010011101;
        a_array[34] = 32'b00111111000000110011010110000101;
        b_array[34] = 32'b00111111001010101110111111110010;
        c_array[34] = 32'b00111111100101110001001010111100;
        a_array[35] = 32'b00111111000010000001011101011100;
        b_array[35] = 32'b00111101001000001110010001101101;
        c_array[35] = 32'b00111111000100100010010110100011;
        a_array[36] = 32'b00111110111000000001001000001001;
        b_array[36] = 32'b00111111011011101000110010111110;
        c_array[36] = 32'b00111111101011110100101011100001;
        a_array[37] = 32'b00111111011011100100100110001101;
        b_array[37] = 32'b00111111001110001001000001010101;
        c_array[37] = 32'b00111111110100110110110011110001;
        a_array[38] = 32'b00111110100100011000111011101000;
        b_array[38] = 32'b00111111001111010001000010010110;
        c_array[38] = 32'b00111111100000101110110000000101;
        a_array[39] = 32'b00111111001000111101010110100111;
        b_array[39] = 32'b00111110101101010100010111011110;
        c_array[39] = 32'b00111111011111100111100010010110;
        a_array[40] = 32'b00111111001100000001011110101111;
        b_array[40] = 32'b00111110001010011111010100100010;
        c_array[40] = 32'b00111111010110101001010011111000;
        a_array[41] = 32'b00111110111000010101010101100001;
        b_array[41] = 32'b00111111011000010100110010011100;
        c_array[41] = 32'b00111111101010001111101110100110;
        a_array[42] = 32'b00111111010101000100011010000110;
        b_array[42] = 32'b00111110101010010010000111110011;
        c_array[42] = 32'b00111111100101000110101111000000;
        a_array[43] = 32'b00111110011010100111011010100010;
        b_array[43] = 32'b00111111011001001011010000001110;
        c_array[43] = 32'b00111111100011111010100011011011;
        a_array[44] = 32'b00111110101100110110001001101001;
        b_array[44] = 32'b00111111001011111100100110011001;
        c_array[44] = 32'b00111111100001001011110101100111;
        a_array[45] = 32'b00111111011101001101101100011010;
        b_array[45] = 32'b00111111000101101011000100011111;
        c_array[45] = 32'b00111111110001011100011000011100;
        a_array[46] = 32'b00111111001010000100010100010100;
        b_array[46] = 32'b00111111010110111101001000110110;
        c_array[46] = 32'b00111111110000100000101110100101;
        a_array[47] = 32'b00111110111000010000110111111111;
        b_array[47] = 32'b00111111011011001000100101001001;
        c_array[47] = 32'b00111111101011101000100000100100;
        a_array[48] = 32'b00111110110010111111111111100100;
        b_array[48] = 32'b00111111010100001001010010010000;
        c_array[48] = 32'b00111111100110110100101001000001;
        a_array[49] = 32'b00111111001011110010100011110010;
        b_array[49] = 32'b00111111011010010011010101110111;
        c_array[49] = 32'b00111111110011000010111100110100;
        a_array[50] = 32'b00111110111101110000100100000100;
        b_array[50] = 32'b00111110010111010000000100111000;
        c_array[50] = 32'b00111111001100101100010011010000;
        a_array[51] = 32'b00111111011100110100001110111101;
        b_array[51] = 32'b00111111011010111000110110000110;
        c_array[51] = 32'b00111111111011110110100010100010;
        a_array[52] = 32'b00111110000101110011010000110000;
        b_array[52] = 32'b00111111011000011000110101001010;
        c_array[52] = 32'b00111111100000111010110100101011;
        a_array[53] = 32'b00111111001001000001110111011100;
        b_array[53] = 32'b00111110110111010010100100000000;
        c_array[53] = 32'b00111111100010010101100100101110;
        a_array[54] = 32'b00111111000111101001110111100000;
        b_array[54] = 32'b00111110100011111110011100000101;
        c_array[54] = 32'b00111111011001101001000101100010;
        a_array[55] = 32'b00111111010010010011011101101111;
        b_array[55] = 32'b00111110100111010110101100011110;
        c_array[55] = 32'b00111111100010111111011001111111;
        a_array[56] = 32'b00111110111001001110000110010110;
        b_array[56] = 32'b00111110011001111000100001111111;
        c_array[56] = 32'b00111111001011000101001011101011;
        a_array[57] = 32'b00111110010000000000100010101110;
        b_array[57] = 32'b00111110100011010110111010100010;
        c_array[57] = 32'b00111110111011010111001011111001;
        a_array[58] = 32'b00111111000011100111001100011001;
        b_array[58] = 32'b00111110110101010011111110101000;
        c_array[58] = 32'b00111111011110010001001011101101;
        a_array[59] = 32'b00111110001011011010110101111011;
        b_array[59] = 32'b00111111011010000010010001001101;
        c_array[59] = 32'b00111111100010011100011111010110;
        a_array[60] = 32'b00111101110100110100101101101010;
        b_array[60] = 32'b00111110000000010001100111100101;
        c_array[60] = 32'b00111110011010101011111110011010;
        a_array[61] = 32'b00111110111111011010101011011000;
        b_array[61] = 32'b00111111010000101010111010000001;
        c_array[61] = 32'b00111111101000001100000111110110;
        a_array[62] = 32'b00111111011111000001100010101111;
        b_array[62] = 32'b00111111011011110101110001101100;
        c_array[62] = 32'b00111111111101011011101010001110;
        a_array[63] = 32'b00111111001011110011011111001010;
        b_array[63] = 32'b00111110110001000011000101000011;
        c_array[63] = 32'b00111111100010001010100000110110;
        a_array[64] = 32'b00111111001111111111000011111100;
        b_array[64] = 32'b00111110101111001100000101111000;
        c_array[64] = 32'b00111111100011110010100011011100;
        a_array[65] = 32'b00111110100101101001110000110000;
        b_array[65] = 32'b00111110011011011101010111111000;
        c_array[65] = 32'b00111111000001101100001110010110;
        a_array[66] = 32'b00111111000101011010000100001010;
        b_array[66] = 32'b00111110011110100100011101010101;
        c_array[66] = 32'b00111111010101000011001011011111;
        a_array[67] = 32'b00111110000111000000110000010010;
        b_array[67] = 32'b00111111001110110110111000010110;
        c_array[67] = 32'b00111111011000100111000100011010;
        a_array[68] = 32'b00111110000000000111110001111110;
        b_array[68] = 32'b00111111010010110010000011100000;
        c_array[68] = 32'b00111111011010110100000000000000;
        a_array[69] = 32'b00111110001010000000101001010110;
        b_array[69] = 32'b00111111001111101011110100000000;
        c_array[69] = 32'b00111111011010001011111110010110;
        a_array[70] = 32'b00111101100110001010001100010100;
        b_array[70] = 32'b00111111011100110011101000000101;
        c_array[70] = 32'b00111111100000110010011100110100;
        a_array[71] = 32'b00111101010101110010100011101100;
        b_array[71] = 32'b00111111000001011000010100101101;
        c_array[71] = 32'b00111111000100101111011110111100;
        a_array[72] = 32'b00111110001101000111000010010001;
        b_array[72] = 32'b00111110011101011101001011101001;
        c_array[72] = 32'b00111110110101010010000110111101;
        a_array[73] = 32'b00111111010011000011110001111110;
        b_array[73] = 32'b00111111001110111000111100111101;
        c_array[73] = 32'b00111111110000111110010111011110;
        a_array[74] = 32'b00111111001010000001010010001110;
        b_array[74] = 32'b00111111011101111010011111011101;
        c_array[74] = 32'b00111111110011111101111000110110;
        a_array[75] = 32'b00111111001000111011001110001011;
        b_array[75] = 32'b00111111010000100111110111111100;
        c_array[75] = 32'b00111111101100110001100011000100;
        a_array[76] = 32'b00111101101111110111001010110001;
        b_array[76] = 32'b00111110000010100010001111011100;
        c_array[76] = 32'b00111110011010011101110100110100;
        a_array[77] = 32'b00111111000001010010110001111101;
        b_array[77] = 32'b00111101101000000011100000101100;
        c_array[77] = 32'b00111111000110010011001110000010;
        a_array[78] = 32'b00111101100011110010101100010110;
        b_array[78] = 32'b00111110010100011001000100011010;
        c_array[78] = 32'b00111110100011001001001101010010;
        a_array[79] = 32'b00111110111011000011111101001110;
        b_array[79] = 32'b00111111010100011101011001011111;
        c_array[79] = 32'b00111111101000111111101100000011;
        a_array[80] = 32'b00111111000100101100010100000010;
        b_array[80] = 32'b00111111010000010110110110111111;
        c_array[80] = 32'b00111111101010100001100101100000;
        a_array[81] = 32'b00111101010101001011110111001100;
        b_array[81] = 32'b00111110001000011001100000110001;
        c_array[81] = 32'b00111110010101101100011110100100;
        a_array[82] = 32'b00111111011111111111111110010100;
        b_array[82] = 32'b00111110010100010011101110000101;
        c_array[82] = 32'b00111111100110100010011100111011;
        a_array[83] = 32'b00111111011000111101010000100010;
        b_array[83] = 32'b00111110000000000111101011001111;
        c_array[83] = 32'b00111111100000011111100101101011;
        a_array[84] = 32'b00111111011111110110111111000001;
        b_array[84] = 32'b00111101010111010110101101111010;
        c_array[84] = 32'b00111111100001101010001100111100;
        a_array[85] = 32'b00111111010111101101101110110011;
        b_array[85] = 32'b00111101100101000010000100011111;
        c_array[85] = 32'b00111111011100010101111111010111;
        a_array[86] = 32'b00111011100010000101111000011011;
        b_array[86] = 32'b00111111011011000100111001000010;
        c_array[86] = 32'b00111111011011010101111011111110;
        a_array[87] = 32'b00111111000110000000100101010001;
        b_array[87] = 32'b00111110001110001011001110000010;
        c_array[87] = 32'b00111111010001100011011000110010;
        a_array[88] = 32'b00111110001001110000101111110010;
        b_array[88] = 32'b00111110110010001000101110011111;
        c_array[88] = 32'b00111111000011100000100011001100;
        a_array[89] = 32'b00111111011010011011110000011110;
        b_array[89] = 32'b00111111010100011101011110001011;
        c_array[89] = 32'b00111111110111011100100111010100;
        a_array[90] = 32'b00111110101101111101101101011001;
        b_array[90] = 32'b00111111000011010110111110101001;
        c_array[90] = 32'b00111111011010010101110101010110;
        a_array[91] = 32'b00111111000101000101010110000110;
        b_array[91] = 32'b00111110111001111011100000000101;
        c_array[91] = 32'b00111111100001000001100011000100;
        a_array[92] = 32'b00111111001011111111100010011111;
        b_array[92] = 32'b00111101110011000001000000010111;
        c_array[92] = 32'b00111111010010010111101010100010;
        a_array[93] = 32'b00111111000001111110001100001000;
        b_array[93] = 32'b00111111010000011101111000000010;
        c_array[93] = 32'b00111111101001001110000010000101;
        a_array[94] = 32'b00111110100110111100110010010011;
        b_array[94] = 32'b00111111011111100000001010101111;
        c_array[94] = 32'b00111111101001011111010001111100;
        a_array[95] = 32'b00111111000100111011010001100001;
        b_array[95] = 32'b00111111011000001010101101001100;
        c_array[95] = 32'b00111111101110100010111111010110;
        a_array[96] = 32'b00111111001111110111000001101110;
        b_array[96] = 32'b00111111001000010000000000111110;
        c_array[96] = 32'b00111111101100000011100001010110;
        a_array[97] = 32'b00111101000100010001010110000011;
        b_array[97] = 32'b00111111001111110111000000000010;
        c_array[97] = 32'b00111111010010001000000101011010;
        a_array[98] = 32'b00111111010101010100111100011111;
        b_array[98] = 32'b00111111011011001110010101111010;
        c_array[98] = 32'b00111111111000010001101001001100;
        a_array[99] = 32'b00111111010111111000111010110110;
        b_array[99] = 32'b00111111010101001011111011100000;
        c_array[99] = 32'b00111111110110100010011011001011;
        for (i = 0; i < 100; i = i + 1) begin
            rst = 0;
            #10;
            rst = 1;
            a = a_array[i];
            b = b_array[i];
            for (j = 0; j < 100; j = j + 1) begin
//                $display("state: %d, c: %b", state, c);
                #10;
            end
            if (c !== c_array[i]) begin
                 $display("Wrong Answer! a: %b, b: %b, output: %b, expected: %b", a, b, c, c_array[i]);
                 $fatal;
            end
        end
		$display("Congratulations! You have passed all of the tests.");
		$finish;
    end
endmodule