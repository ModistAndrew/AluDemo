`include "float_adder.v"

module test_float_adder;
    reg clk = 1;
    always #5 clk = ~clk;
    reg [31:0] a, b;
    wire [31:0] c;
    wire [2:0] state;
    reg rst;
    reg [31:0] a_array [0:99];
    reg [31:0] b_array [0:99];
    reg [31:0] c_array [0:99];
    FAdd float_adder(
        .clk(clk),
        .rst(rst),
        .a(a),
        .b(b),
        .c(c),
        .state(state)
    );
    integer i;
    integer j;
    initial begin

a_array[0] = 32'b01101011100010110100010101100111;
b_array[0] = 32'b11100100001111001001100001101001;
c_array[0] = 32'b01101011100010110100001111101110;
a_array[1] = 32'b11110100101100001101110001010001;
b_array[1] = 32'b00101010111010001001010001001010;
c_array[1] = 32'b11110100101100001101110001010001;
a_array[2] = 32'b10100011100011100001111100101001;
b_array[2] = 32'b10111101000110110101100010111010;
c_array[2] = 32'b10111101000110110101100010111010;
a_array[3] = 32'b10101110101100010100000111110010;
b_array[3] = 32'b01111001111000101010100111100011;
c_array[3] = 32'b01111001111000101010100111100011;
a_array[4] = 32'b01010001010111110000000001111100;
b_array[4] = 32'b00010010001000000000100001010100;
c_array[4] = 32'b01010001010111110000000001111100;
a_array[5] = 32'b00000010000101100010001100011011;
b_array[5] = 32'b10010001100100001100110111100111;
c_array[5] = 32'b10010001100100001100110111100111;
a_array[6] = 32'b00010100000011100000111101110110;
b_array[6] = 32'b10010000100111001111100100101110;
c_array[6] = 32'b00010100000011001101010110000100;
a_array[7] = 32'b11111111110111001100001000110011;
b_array[7] = 32'b01000001101001111100010011001001;
c_array[7] = 32'b11111111110111001100001000110011;
a_array[8] = 32'b01001110011010101111101101100110;
b_array[8] = 32'b11010001100110110101000000001101;
c_array[8] = 32'b11010001100110010111101000010110;
a_array[9] = 32'b00111111001011011011101000110001;
b_array[9] = 32'b00100101011100010011000010100011;
c_array[9] = 32'b00111111001011011011101000110001;
a_array[10] = 32'b11000011011011000110000100100101;
b_array[10] = 32'b10110011001110101011000100000101;
c_array[10] = 32'b11000011011011000110000100100101;
a_array[11] = 32'b10100100010000111010100001011000;
b_array[11] = 32'b01100111011000111000010001011110;
c_array[11] = 32'b01100111011000111000010001011110;
a_array[12] = 32'b00001000111011011011110110101011;
b_array[12] = 32'b01000011010100111101000011001101;
c_array[12] = 32'b01000011010100111101000011001101;
a_array[13] = 32'b00011000100110100111011010011011;
b_array[13] = 32'b11110001111100110010010001010100;
c_array[13] = 32'b11110001111100110010010001010100;
a_array[14] = 32'b00001000001101101100010000001110;
b_array[14] = 32'b10111010100101011111100001110100;
c_array[14] = 32'b10111010100101011111100001110100;
a_array[15] = 32'b10011110011111111111010100100001;
b_array[15] = 32'b11110011011110111000110111011100;
c_array[15] = 32'b11110011011110111000110111011100;
a_array[16] = 32'b10100010001000100001101001110000;
b_array[16] = 32'b10110000000001101100100000111110;
c_array[16] = 32'b10110000000001101100100000111110;
a_array[17] = 32'b11000001100110101100001001000001;
b_array[17] = 32'b11000100000010111010110111111100;
c_array[17] = 32'b11000100000100001000010000001110;
a_array[18] = 32'b10111000000001001000001000111110;
b_array[18] = 32'b11110111001001001100011001111110;
c_array[18] = 32'b11110111001001001100011001111110;
a_array[19] = 32'b00100100011000111011100111101010;
b_array[19] = 32'b01010001111010101101001101101011;
c_array[19] = 32'b01010001111010101101001101101011;
a_array[20] = 32'b01011000000010111101011110001111;
b_array[20] = 32'b00111000010101010101100001011100;
c_array[20] = 32'b01011000000010111101011110001111;
a_array[21] = 32'b01101010001000110100001011101100;
b_array[21] = 32'b10011101010011101101010000111011;
c_array[21] = 32'b01101010001000110100001011101100;
a_array[22] = 32'b10101100110110001001101000110010;
b_array[22] = 32'b01111010011011011000110100111100;
c_array[22] = 32'b01111010011011011000110100111100;
a_array[23] = 32'b01010100001000101000100111101100;
b_array[23] = 32'b00111000010000110111111111011011;
c_array[23] = 32'b01010100001000101000100111101100;
a_array[24] = 32'b00110010111111111111100100000010;
b_array[24] = 32'b11010111100101000111100011111110;
c_array[24] = 32'b11010111100101000111100011111110;
a_array[25] = 32'b00111101110000100100000011111011;
b_array[25] = 32'b01111001101000011101111010101010;
c_array[25] = 32'b01111001101000011101111010101010;
a_array[26] = 32'b10010010111001101000010111111011;
b_array[26] = 32'b01010010000011101110110111010001;
c_array[26] = 32'b01010010000011101110110111010001;
a_array[27] = 32'b01001111010011101111000000000101;
b_array[27] = 32'b01100100100110111011011101111100;
c_array[27] = 32'b01100100100110111011011101111100;
a_array[28] = 32'b00111001001110000110010101110101;
b_array[28] = 32'b10011000000000010001010110111110;
c_array[28] = 32'b00111001001110000110010101110101;
a_array[29] = 32'b11000111001110011000110010001001;
b_array[29] = 32'b10010101101101011010111101011100;
c_array[29] = 32'b11000111001110011000110010001001;
a_array[30] = 32'b10001101001101001011011010101000;
b_array[30] = 32'b10111111011010101011011000001111;
c_array[30] = 32'b10111111011010101011011000001111;
a_array[31] = 32'b11111110000011000101011110110001;
b_array[31] = 32'b11010111100110111110010011110001;
c_array[31] = 32'b11111110000011000101011110110001;
a_array[32] = 32'b11011111111110000111111000000101;
b_array[32] = 32'b00100101101001110000101111110111;
c_array[32] = 32'b11011111111110000111111000000101;
a_array[33] = 32'b11001010110100001000010011101001;
b_array[33] = 32'b10010011100000011000001000111010;
c_array[33] = 32'b11001010110100001000010011101001;
a_array[34] = 32'b10010000000011111000111111001010;
b_array[34] = 32'b00010101000000010100101011001011;
c_array[34] = 32'b00010101000000010010011011100111;
a_array[35] = 32'b10001001100010100011000101001000;
b_array[35] = 32'b10000110101110010100011101100100;
c_array[35] = 32'b10001001100011010001011001100110;
a_array[36] = 32'b10010110100011100001001000011111;
b_array[36] = 32'b01100110000111100011111100011110;
c_array[36] = 32'b01100110000111100011111100011110;
a_array[37] = 32'b11010100000010100100011100011100;
b_array[37] = 32'b11010001110110011100010101100100;
c_array[37] = 32'b11010100000100010001010101000111;
a_array[38] = 32'b10001011111101110010101100010100;
b_array[38] = 32'b11000010100101100011111001011010;
c_array[38] = 32'b11000010100101100011111001011010;
a_array[39] = 32'b10001000111100101011000101011110;
b_array[39] = 32'b10111011000011111101001101111001;
c_array[39] = 32'b10111011000011111101001101111001;
a_array[40] = 32'b01001001011000101000000100111011;
b_array[40] = 32'b00000110101001011110111001100100;
c_array[40] = 32'b01001001011000101000000100111011;
a_array[41] = 32'b01111111111111111100101000010001;
b_array[41] = 32'b01110001111010100001000100001001;
c_array[41] = 32'b01111111111111111100101000010001;
a_array[42] = 32'b01111111101101111110000010101010;
b_array[42] = 32'b01101111011011011101100110101100;
c_array[42] = 32'b01111111111101111110000010101010;
a_array[43] = 32'b00000000100010000101111000011011;
b_array[43] = 32'b11001100000001001010100010101111;
c_array[43] = 32'b11001100000001001010100010101111;
a_array[44] = 32'b10010100111000010111111000110011;
b_array[44] = 32'b01110100110111100000111011100011;
c_array[44] = 32'b01110100110111100000111011100011;
a_array[45] = 32'b10101101111101101101011001001000;
b_array[45] = 32'b01001010001010101100001100010101;
c_array[45] = 32'b01001010001010101100001100010101;
a_array[46] = 32'b11010111111111000100111110111011;
b_array[46] = 32'b11000011111100011000010000100010;
c_array[46] = 32'b11010111111111000100111110111011;
a_array[47] = 32'b10100110111100110010010010111010;
b_array[47] = 32'b11001001110110100011000001111101;
c_array[47] = 32'b11001001110110100011000001111101;
a_array[48] = 32'b11011111101110000011011100001011;
b_array[48] = 32'b00000100100010001010110000011010;
c_array[48] = 32'b11011111101110000011011100001011;
a_array[49] = 32'b11101010101001111000111101111111;
b_array[49] = 32'b11101111110001110101101011111000;
c_array[49] = 32'b11101111110001111000010011011100;
a_array[50] = 32'b01111101010111100001100011111000;
b_array[50] = 32'b11110011101000011000001000011011;
c_array[50] = 32'b01111101010111100001100011100100;
a_array[51] = 32'b01010101010111000101010110110101;
b_array[51] = 32'b00010100111111001110011101001110;
c_array[51] = 32'b01010101010111000101010110110101;
a_array[52] = 32'b01110001110010010001001010011000;
b_array[52] = 32'b01010011001010011001100100111000;
c_array[52] = 32'b01110001110010010001001010011000;
a_array[53] = 32'b11010000100100101100101001111001;
b_array[53] = 32'b01011001101011011110101000111101;
c_array[53] = 32'b01011001101011011110101000011000;
a_array[54] = 32'b10101010000101010101110110111100;
b_array[54] = 32'b10001001011111100001101101001110;
c_array[54] = 32'b10101010000101010101110110111100;
a_array[55] = 32'b10011100101000001100010111111010;
b_array[55] = 32'b11000001010111100010100001101100;
c_array[55] = 32'b11000001010111100010100001101100;
a_array[56] = 32'b00100011110110000110101010101100;
b_array[56] = 32'b11011100000100001111111000100001;
c_array[56] = 32'b11011100000100001111111000100001;
a_array[57] = 32'b00111100010110011001000110101010;
b_array[57] = 32'b01111000110111110110101001010101;
c_array[57] = 32'b01111000110111110110101001010101;
a_array[58] = 32'b00101011000011011000110110111110;
b_array[58] = 32'b10110111100111100010000110110101;
c_array[58] = 32'b10110111100111100010000110110101;
a_array[59] = 32'b00101100001001110001011100111011;
b_array[59] = 32'b11101010101001111011011101011100;
c_array[59] = 32'b11101010101001111011011101011100;
a_array[60] = 32'b01010110011101011111111100110110;
b_array[60] = 32'b10111101101100000001001010110011;
c_array[60] = 32'b01010110011101011111111100110110;
a_array[61] = 32'b01011011001001011010110011100010;
b_array[61] = 32'b01001111100101111110001111100100;
c_array[61] = 32'b01011011001001011010110011100011;
a_array[62] = 32'b00110100111111010110101101001111;
b_array[62] = 32'b11010110010000111000110100010101;
c_array[62] = 32'b11010110010000111000110100010101;
a_array[63] = 32'b00101100011011100100101011111101;
b_array[63] = 32'b11001101111101110010111001001110;
c_array[63] = 32'b11001101111101110010111001001110;
a_array[64] = 32'b01011101100010001000101000001000;
b_array[64] = 32'b01011110110001101010111111010100;
c_array[64] = 32'b01011110111010001101001001010110;
a_array[65] = 32'b11110101111000001000010110001010;
b_array[65] = 32'b01010011100110011100011001010100;
c_array[65] = 32'b11110101111000001000010110001010;
a_array[66] = 32'b01000100001001110000011010011010;
b_array[66] = 32'b10100001010101111111011010111100;
c_array[66] = 32'b01000100001001110000011010011010;
a_array[67] = 32'b01010111110100101111000100001110;
b_array[67] = 32'b00001110001111100100011110101000;
c_array[67] = 32'b01010111110100101111000100001110;
a_array[68] = 32'b11001001110100001111111010101100;
b_array[68] = 32'b01010101010100011011100111110011;
c_array[68] = 32'b01010101010100011011100111110001;
a_array[69] = 32'b11100011010011000101011101001100;
b_array[69] = 32'b10101010001100011011011000101101;
c_array[69] = 32'b11100011010011000101011101001100;
a_array[70] = 32'b01111101111111111001110100001001;
b_array[70] = 32'b01101001111001111111001111100101;
c_array[70] = 32'b01111101111111111001110100001001;
a_array[71] = 32'b10011000000101101111100011000100;
b_array[71] = 32'b11111010101101001001110110101111;
c_array[71] = 32'b11111010101101001001110110101111;
a_array[72] = 32'b01100001111001110100111010100011;
b_array[72] = 32'b10001111100000011001111001111111;
c_array[72] = 32'b01100001111001110100111010100011;
a_array[73] = 32'b00110001001000010110011110101101;
b_array[73] = 32'b11111000101101011110011101110110;
c_array[73] = 32'b11111000101101011110011101110110;
a_array[74] = 32'b01101110010100110100110011011110;
b_array[74] = 32'b01100101100101101000110000011100;
c_array[74] = 32'b01101110010100110100110100101001;
a_array[75] = 32'b00100110000011011000110001001010;
b_array[75] = 32'b01110100011011110010111000110000;
c_array[75] = 32'b01110100011011110010111000110000;
a_array[76] = 32'b10111111110000110010111000100000;
b_array[76] = 32'b00010100110101010011011010000101;
c_array[76] = 32'b10111111110000110010111000100000;
a_array[77] = 32'b01101110101010101000010111111011;
b_array[77] = 32'b00111011010110010100100000000111;
c_array[77] = 32'b01101110101010101000010111111011;
a_array[78] = 32'b00111111011111000010111111110100;
b_array[78] = 32'b10010111000110000000101100001011;
c_array[78] = 32'b00111111011111000010111111110100;
a_array[79] = 32'b01011101001000000101111000100000;
b_array[79] = 32'b11001101001100101010101110000110;
c_array[79] = 32'b01011101001000000101111000100000;
a_array[80] = 32'b11101011010001111111011000111110;
b_array[80] = 32'b00010110110011111000000011110001;
c_array[80] = 32'b11101011010001111111011000111110;
a_array[81] = 32'b10111111110011111010111011011001;
b_array[81] = 32'b10010001101100011100110000110011;
c_array[81] = 32'b10111111110011111010111011011001;
a_array[82] = 32'b00101001100100110100011010011001;
b_array[82] = 32'b11110100010010010011100110100011;
c_array[82] = 32'b11110100010010010011100110100011;
a_array[83] = 32'b11101011000111010010110000010100;
b_array[83] = 32'b00111111011111110101110111011001;
c_array[83] = 32'b11101011000111010010110000010100;
a_array[84] = 32'b00110010011110010100111111110111;
b_array[84] = 32'b01001101111011111101111110100000;
c_array[84] = 32'b01001101111011111101111110100000;
a_array[85] = 32'b00010011010110111000000100010000;
b_array[85] = 32'b10001101110011011111100011110110;
c_array[85] = 32'b00010011010110110110011101010001;
a_array[86] = 32'b10101110100010100110001110010100;
b_array[86] = 32'b00101010011010101101100110111110;
c_array[86] = 32'b10101110100010011110111000100111;
a_array[87] = 32'b00110110101100101010110010111100;
b_array[87] = 32'b01001010101100100110111001111000;
c_array[87] = 32'b01001010101100100110111001111000;
a_array[88] = 32'b11010100010100011100111101001001;
b_array[88] = 32'b10111110011001000000000011100110;
c_array[88] = 32'b11010100010100011100111101001001;
a_array[89] = 32'b01110001000001110101011111010000;
b_array[89] = 32'b11000010010001000111100111011010;
c_array[89] = 32'b01110001000001110101011111010000;
a_array[90] = 32'b01000111010111100010010101101010;
b_array[90] = 32'b01101010001110110111000101001100;
c_array[90] = 32'b01101010001110110111000101001100;
a_array[91] = 32'b10011111010001100001101101010001;
b_array[91] = 32'b01011101010110111010101110110011;
c_array[91] = 32'b01011101010110111010101110110011;
a_array[92] = 32'b11111110000011110110001110000100;
b_array[92] = 32'b01110010111000110100000100111010;
c_array[92] = 32'b11111110000011110110001110000010;
a_array[93] = 32'b10110100100101001011001011111011;
b_array[93] = 32'b01100100010000101001010110011001;
c_array[93] = 32'b01100100010000101001010110011001;
a_array[94] = 32'b10100101100101110011111000110010;
b_array[94] = 32'b01101110110010011101100001000100;
c_array[94] = 32'b01101110110010011101100001000100;
a_array[95] = 32'b00000110010010101111010010011011;
b_array[95] = 32'b11111110010001001000110111101001;
c_array[95] = 32'b11111110010001001000110111101001;
a_array[96] = 32'b10011010111111100011011000100101;
b_array[96] = 32'b11101110101111100100001000001000;
c_array[96] = 32'b11101110101111100100001000001000;
a_array[97] = 32'b00001100101111100101101111101001;
b_array[97] = 32'b10100110101000000010110001011110;
c_array[97] = 32'b10100110101000000010110001011110;
a_array[98] = 32'b01100111100100000110111101100000;
b_array[98] = 32'b00000110100101111101001011010010;
c_array[98] = 32'b01100111100100000110111101100000;
a_array[99] = 32'b10111010100101100110110011010000;
b_array[99] = 32'b01011000100101011111010111111010;
c_array[99] = 32'b01011000100101011111010111111010;
        #5;
        for (i = 0; i < 100; i = i + 1) begin
            rst = 0;
            #10;
            rst = 1;
            a = a_array[i];
            b = b_array[i];
            for (j = 0; j < 300; j = j + 1) begin // it takes at most about 255 + 32 cycles to finish the calculation
//                $display("state: %d, c: %b", state, c);
                #10;
            end
            if (c !== c_array[i] && !(c === 32'b01111111100000000000000000000001 && c_array[i][30:23] === 8'b11111111 && c_array[i][22:0] !== 23'b0)) begin
                 $display("Wrong Answer! i: %d, a: %b, b: %b, output: %b, expected: %b", i, a, b, c, c_array[i]);
                 $fatal;
            end
        end
		$display("Congratulations! You have passed all of the tests.");
		$finish;
    end
endmodule